`timescale 1ns / 1ps

module dithering(

    );
    
    
endmodule
